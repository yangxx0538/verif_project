/*

Copyright (c) 2014-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * Priority encoder module
 */
module verif_priority_encoder #
(
    parameter WIDTH = 4,
    // LSB priority: "LOW", "HIGH"
    parameter LSB_PRIORITY = "LOW"
)
(
    input wire [WIDTH-1:0]         input_unencoded,
    input wire                     output_valid,
    input wire [$clog2(WIDTH)-1:0] output_encoded,
    input wire [WIDTH-1:0]         output_unencoded
);

assert property (
	output_valid & (!input_unencoded[0] &!input_unencoded[1])
);

endmodule


module Wrapper;

bind priority_encoder verif_priority_encoder # ( 
		.WIDTH(WIDTH),
		.LSB_PRIORITY(LSB_PRIORITY)
		
	) verif_priority_encoder_inst (
		.input_unencoded(input_unencoded),
		.output_valid(output_valid),
		.output_encoded(output_encoded),
		.output_unencoded(output_unencoded)
	);

endmodule